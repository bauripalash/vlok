module lib

//Transaction structure of block data
pub struct Transaction {
pub mut:
	from   string
	to     string
	amount u64
}
