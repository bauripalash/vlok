module lib

// TODO: Blockchain server
